library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity somador is
PORT(
		entradaA : in 	std_logic_vector(15 downto 0);
		entradaB : in 	std_logic_vector(15 downto 0);
		saida 	: out std_logic_vector(15 downto 0));
end somador;
	
architecture hardware of somador is

	signal entrada_A 	: std_logic_vector(15 downto 0);
	signal entrada_B 	: std_logic_vector(15 downto 0);
	signal saida_soma : std_logic_vector(15 downto 0);

	component somador_16bits
		PORT(
			entradaA : in 	std_logic_vector(15 downto 0);
			entradaB : in 	std_logic_vector(15 downto 0);
			saida 	: out std_logic_vector(15 downto 0));
	end component;

begin

	saida_soma(15 downto 0) <= ("0000000000000000" & entradaA(15 downto 0)) + ("0000000000000000" & entradaB(15 downto 0));
	
	rot_soma : somador_16bits PORT MAP
	(
		entradaA => entrada_A,
		entradaB => entrada_B,
		saida 	=> saida_soma	
	);
	
	signal_a_somador : process
	begin
		entrada_A <= "0000000000000000"; wait for 50 ns;
		entrada_A <= "0000000000000001"; wait for 50 ns;
		entrada_A <= "0000000000000010"; wait for 50 ns;
		entrada_A <= "0000000000000011"; wait for 50 ns;
		entrada_A <= "0000000000000100"; wait for 50 ns;
		entrada_A <= "0000000000000101"; wait for 50 ns;
		entrada_A <= "0000000000000110"; wait for 50 ns;
		entrada_A <= "0000000000000111"; wait for 50 ns;
		entrada_A <= "0000000000001000"; wait for 50 ns;
		entrada_A <= "0000000000001001"; wait for 50 ns;
		entrada_A <= "0000000000001010"; wait for 50 ns;
		entrada_A <= "0000000000001011"; wait for 50 ns;
		entrada_A <= "0000000000001100"; wait for 50 ns;
		entrada_A <= "0000000000001101"; wait for 50 ns;
		entrada_A <= "0000000000001111"; wait for 50 ns;
		entrada_A <= "0000000000010000"; wait for 50 ns;
		entrada_A <= "0000000000010001"; wait for 50 ns;
		entrada_A <= "0000000000010010"; wait for 50 ns;
		entrada_A <= "0000000000010011"; wait for 50 ns;
		entrada_A <= "0000000000010100"; wait for 50 ns;
		entrada_A <= "0000000000010101"; wait for 50 ns;
		entrada_A <= "0000000000010110"; wait for 50 ns;
		entrada_A <= "0000000000010111"; wait for 50 ns;
		entrada_A <= "0000000000011000"; wait for 50 ns;
		entrada_A <= "0000000000011001"; wait for 50 ns;
		entrada_A <= "0000000000011010"; wait for 50 ns;
		entrada_A <= "0000000000011011"; wait for 50 ns;
		entrada_A <= "0000000000011100"; wait for 50 ns;
		entrada_A <= "0000000000011101"; wait for 50 ns;
		entrada_A <= "0000000000011110"; wait for 50 ns;
		entrada_A <= "0000000000011111"; wait for 50 ns;
		entrada_A <= "0000000000100000"; wait for 50 ns;
		entrada_A <= "0000000000100001"; wait for 50 ns;
		entrada_A <= "0000000000100010"; wait for 50 ns;
		entrada_A <= "0000000000100011"; wait for 50 ns;
		entrada_A <= "0000000000100100"; wait for 50 ns;
		entrada_A <= "0000000000100101"; wait for 50 ns;
		entrada_A <= "0000000000100110"; wait for 50 ns;
		entrada_A <= "0000000000100111"; wait for 50 ns;
		entrada_A <= "0000000000101000"; wait for 50 ns;
		entrada_A <= "0000000000101001"; wait for 50 ns;
		entrada_A <= "0000000000101010"; wait for 50 ns;
		entrada_A <= "0000000000101011"; wait for 50 ns;
		entrada_A <= "0000000000101100"; wait for 50 ns;
		entrada_A <= "0000000000101101"; wait for 50 ns;
		entrada_A <= "0000000000101110"; wait for 50 ns;
		entrada_A <= "0000000000101111"; wait for 50 ns;
		entrada_A <= "0000000000110000"; wait for 50 ns;
		entrada_A <= "0000000000110001"; wait for 50 ns;
		entrada_A <= "0000000000110010"; wait for 50 ns;
		entrada_A <= "0000000000110011"; wait for 50 ns;
		entrada_A <= "0000000000110100"; wait for 50 ns;
		entrada_A <= "0000000000110101"; wait for 50 ns;
		entrada_A <= "0000000000110110"; wait for 50 ns;
		entrada_A <= "0000000000110111"; wait for 50 ns;
		entrada_A <= "0000000000111000"; wait for 50 ns;
		entrada_A <= "0000000000111001"; wait for 50 ns;
		entrada_A <= "0000000000111010"; wait for 50 ns;
		entrada_A <= "0000000000111011"; wait for 50 ns;
		entrada_A <= "0000000000111100"; wait for 50 ns;
		entrada_A <= "0000000000111101"; wait for 50 ns;
		entrada_A <= "0000000000111110"; wait for 50 ns;
		entrada_A <= "0000000000111111"; wait for 50 ns;
		entrada_A <= "0000000001000000"; wait for 50 ns;
		entrada_A <= "0000000001000001"; wait for 50 ns;
		entrada_A <= "0000000001000010"; wait for 50 ns;
		entrada_A <= "0000000001000011"; wait for 50 ns;
		entrada_A <= "0000000001000100"; wait for 50 ns;
		entrada_A <= "0000000001000101"; wait for 50 ns;
		entrada_A <= "0000000001000110"; wait for 50 ns;
		entrada_A <= "0000000001000111"; wait for 50 ns;
		entrada_A <= "0000000001001000"; wait for 50 ns;
		entrada_A <= "0000000001001001"; wait for 50 ns;
		entrada_A <= "0000000001001010"; wait for 50 ns;
		entrada_A <= "0000000001001011"; wait for 50 ns;
		entrada_A <= "0000000001001100"; wait for 50 ns;
		entrada_A <= "0000000001001101"; wait for 50 ns;
		entrada_A <= "0000000001001110"; wait for 50 ns;
		entrada_A <= "0000000001001111"; wait for 50 ns;
		entrada_A <= "0000000001010000"; wait for 50 ns;
		entrada_A <= "0000000001010001"; wait for 50 ns;
		entrada_A <= "0000000001010010"; wait for 50 ns;
		entrada_A <= "0000000001010011"; wait for 50 ns;
		entrada_A <= "0000000001010100"; wait for 50 ns;
		entrada_A <= "0000000001010101"; wait for 50 ns;
		entrada_A <= "0000000001010110"; wait for 50 ns;
		entrada_A <= "0000000001010111"; wait for 50 ns;
		entrada_A <= "0000000001011000"; wait for 50 ns;
		entrada_A <= "0000000001011001"; wait for 50 ns;
		entrada_A <= "0000000001011010"; wait for 50 ns;
		entrada_A <= "0000000001011011"; wait for 50 ns;
		entrada_A <= "0000000001011100"; wait for 50 ns;
		entrada_A <= "0000000001011101"; wait for 50 ns;
		entrada_A <= "0000000001011110"; wait for 50 ns;
		entrada_A <= "0000000001011111"; wait for 50 ns;
		entrada_A <= "0000000001100000"; wait for 50 ns;
		entrada_A <= "0000000001100001"; wait for 50 ns;
		entrada_A <= "0000000001100010"; wait for 50 ns;
		entrada_A <= "0000000001100011"; wait for 50 ns;
		entrada_A <= "0000000001100100"; wait for 50 ns;
		entrada_A <= "0000000001100101"; wait for 50 ns;
		entrada_A <= "0000000001100110"; wait for 50 ns;
		entrada_A <= "0000000001100111"; wait for 50 ns;
		entrada_A <= "0000000001101000"; wait for 50 ns;
		entrada_A <= "0000000001101001"; wait for 50 ns;
		entrada_A <= "0000000001101010"; wait for 50 ns;
		entrada_A <= "0000000001101011"; wait for 50 ns;
		entrada_A <= "0000000001101100"; wait for 50 ns;
		entrada_A <= "0000000001101101"; wait for 50 ns;
		entrada_A <= "0000000001101110"; wait for 50 ns;
		entrada_A <= "0000000001101111"; wait for 50 ns;
		entrada_A <= "0000000001110000"; wait for 50 ns;
		entrada_A <= "0000000001110001"; wait for 50 ns;
		entrada_A <= "0000000001110010"; wait for 50 ns;
		entrada_A <= "0000000001110011"; wait for 50 ns;
		entrada_A <= "0000000001110100"; wait for 50 ns;
		entrada_A <= "0000000001110101"; wait for 50 ns;
		entrada_A <= "0000000001110110"; wait for 50 ns;
		entrada_A <= "0000000001110111"; wait for 50 ns;
		entrada_A <= "0000000001111000"; wait for 50 ns;
		entrada_A <= "0000000001111001"; wait for 50 ns;
		entrada_A <= "0000000001111010"; wait for 50 ns;
		entrada_A <= "0000000001111011"; wait for 50 ns;
		entrada_A <= "0000000001111100"; wait for 50 ns;
		entrada_A <= "0000000001111101"; wait for 50 ns;
		entrada_A <= "0000000001111110"; wait for 50 ns;
		entrada_A <= "0000000001111111"; wait for 50 ns;
		entrada_A <= "0000000010000000"; wait for 50 ns;
		entrada_A <= "0000000010000001"; wait for 50 ns;
		entrada_A <= "0000000010000010"; wait for 50 ns;
		entrada_A <= "0000000010000011"; wait for 50 ns;
		entrada_A <= "0000000010000100"; wait for 50 ns;
		entrada_A <= "0000000010000101"; wait for 50 ns;
		entrada_A <= "0000000010000110"; wait for 50 ns;
		entrada_A <= "0000000010000111"; wait for 50 ns;
		entrada_A <= "0000000010001000"; wait for 50 ns;
		entrada_A <= "0000000010001001"; wait for 50 ns;
		entrada_A <= "0000000010001010"; wait for 50 ns;
		entrada_A <= "0000000010001011"; wait for 50 ns;
		entrada_A <= "0000000010001100"; wait for 50 ns;
		entrada_A <= "0000000010001101"; wait for 50 ns;
		entrada_A <= "0000000010001110"; wait for 50 ns;
		entrada_A <= "0000000010001111"; wait for 50 ns;
		entrada_A <= "0000000010010000"; wait for 50 ns;
		entrada_A <= "0000000010010001"; wait for 50 ns;
		entrada_A <= "0000000010010010"; wait for 50 ns;
		entrada_A <= "0000000010010011"; wait for 50 ns;
		entrada_A <= "0000000010010100"; wait for 50 ns;
		entrada_A <= "0000000010010101"; wait for 50 ns;
		entrada_A <= "0000000010010110"; wait for 50 ns;
		entrada_A <= "0000000010010111"; wait for 50 ns;
		entrada_A <= "0000000010011000"; wait for 50 ns;
		entrada_A <= "0000000010011001"; wait for 50 ns;
		entrada_A <= "0000000010011010"; wait for 50 ns;
		entrada_A <= "0000000010011011"; wait for 50 ns;
		entrada_A <= "0000000010011100"; wait for 50 ns;
		entrada_A <= "0000000010011101"; wait for 50 ns;
		entrada_A <= "0000000010011110"; wait for 50 ns;
		entrada_A <= "0000000010011111"; wait for 50 ns;
		entrada_A <= "0000000010100000"; wait for 50 ns;
		entrada_A <= "0000000010100001"; wait for 50 ns;
		entrada_A <= "0000000010100010"; wait for 50 ns;
		entrada_A <= "0000000010100011"; wait for 50 ns;
		entrada_A <= "0000000010100100"; wait for 50 ns;
		entrada_A <= "0000000010100101"; wait for 50 ns;
		entrada_A <= "0000000010100110"; wait for 50 ns;
		entrada_A <= "0000000010100111"; wait for 50 ns;
		entrada_A <= "0000000010101000"; wait for 50 ns;
		entrada_A <= "0000000010010011"; wait for 50 ns;
		entrada_A <= "0000000010010100"; wait for 50 ns;
		entrada_A <= "0000000010010101"; wait for 50 ns;
		entrada_A <= "0000000010010110"; wait for 50 ns;
		entrada_A <= "0000000010010111"; wait for 50 ns;
		entrada_A <= "0000000010011000"; wait for 50 ns;
		entrada_A <= "0000000010011001"; wait for 50 ns;
		entrada_A <= "0000000010011010"; wait for 50 ns;
		entrada_A <= "0000000010011011"; wait for 50 ns;
		entrada_A <= "0000000010011100"; wait for 50 ns;
		entrada_A <= "0000000010011101"; wait for 50 ns;
		entrada_A <= "0000000010011110"; wait for 50 ns;
		entrada_A <= "0000000010011111"; wait for 50 ns;
		entrada_A <= "0000000010100000"; wait for 50 ns;
		entrada_A <= "0000000010100001"; wait for 50 ns;
		entrada_A <= "0000000010100010"; wait for 50 ns;
		entrada_A <= "0000000010100011"; wait for 50 ns;
		entrada_A <= "0000000010100100"; wait for 50 ns;
		entrada_A <= "0000000010100101"; wait for 50 ns;
		entrada_A <= "0000000010100110"; wait for 50 ns;
		entrada_A <= "0000000010100111"; wait for 50 ns;
		entrada_A <= "0000000010101000"; wait for 50 ns;
		entrada_A <= "0000000010101001"; wait for 50 ns;
		entrada_A <= "0000000010101010"; wait for 50 ns;
		entrada_A <= "0000000010101100"; wait for 50 ns;
		entrada_A <= "0000000010101101"; wait for 50 ns;
		entrada_A <= "0000000010101110"; wait for 50 ns;
		entrada_A <= "0000000010101111"; wait for 50 ns;
		entrada_A <= "0000000010110000"; wait for 50 ns;
		entrada_A <= "0000000010110001"; wait for 50 ns;
		entrada_A <= "0000000010110010"; wait for 50 ns;
		entrada_A <= "0000000010110011"; wait for 50 ns;
		entrada_A <= "0000000010110100"; wait for 50 ns;
		entrada_A <= "0000000010110101"; wait for 50 ns;
		entrada_A <= "0000000010110110"; wait for 50 ns;
		entrada_A <= "0000000010110111"; wait for 50 ns;
		entrada_A <= "0000000010111000"; wait for 50 ns;
		entrada_A <= "0000000010111001"; wait for 50 ns;
		entrada_A <= "0000000010111010"; wait for 50 ns;
		entrada_A <= "0000000010111011"; wait for 50 ns;
		entrada_A <= "0000000010111100"; wait for 50 ns;
		entrada_A <= "0000000010111101"; wait for 50 ns;
		entrada_A <= "0000000010111110"; wait for 50 ns;
		entrada_A <= "0000000010111111"; wait for 50 ns;
		entrada_A <= "0000000011000000"; wait for 50 ns;
		entrada_A <= "0000000011000001"; wait for 50 ns;
		entrada_A <= "0000000011000010"; wait for 50 ns;
		entrada_A <= "0000000011000011"; wait for 50 ns;
		entrada_A <= "0000000011000100"; wait for 50 ns;
		entrada_A <= "0000000011000101"; wait for 50 ns;
		entrada_A <= "0000000011000110"; wait for 50 ns;
		entrada_A <= "0000000011000111"; wait for 50 ns;
		entrada_A <= "0000000011001000"; wait for 50 ns;
		entrada_A <= "0000000011001001"; wait for 50 ns;
		entrada_A <= "0000000011001010"; wait for 50 ns;
		entrada_A <= "0000000011001011"; wait for 50 ns;
		entrada_A <= "0000000011001100"; wait for 50 ns;
		entrada_A <= "0000000011001101"; wait for 50 ns;
		entrada_A <= "0000000011001110"; wait for 50 ns;
		entrada_A <= "0000000011001111"; wait for 50 ns;
		entrada_A <= "0000000011010000"; wait for 50 ns;
		entrada_A <= "0000000011010001"; wait for 50 ns;
		entrada_A <= "0000000011010010"; wait for 50 ns;
		entrada_A <= "0000000011010011"; wait for 50 ns;
		entrada_A <= "0000000011010100"; wait for 50 ns;
		entrada_A <= "0000000011010101"; wait for 50 ns;
		entrada_A <= "0000000011010110"; wait for 50 ns;
		entrada_A <= "0000000011010111"; wait for 50 ns;
		entrada_A <= "0000000011011000"; wait for 50 ns;
		entrada_A <= "0000000011011001"; wait for 50 ns;
		entrada_A <= "0000000011011010"; wait for 50 ns;
		entrada_A <= "0000000011011011"; wait for 50 ns;
		entrada_A <= "0000000011011100"; wait for 50 ns;
		entrada_A <= "0000000011011101"; wait for 50 ns;
		entrada_A <= "0000000011011110"; wait for 50 ns;
		entrada_A <= "0000000011011111"; wait for 50 ns;
		entrada_A <= "0000000011100000"; wait for 50 ns;
		entrada_A <= "0000000011100001"; wait for 50 ns;
		entrada_A <= "0000000011100010"; wait for 50 ns;
		entrada_A <= "0000000011100011"; wait for 50 ns;
		entrada_A <= "0000000011100100"; wait for 50 ns;
		entrada_A <= "0000000011100101"; wait for 50 ns;
		entrada_A <= "0000000011100110"; wait for 50 ns;
		entrada_A <= "0000000011100111"; wait for 50 ns;
		entrada_A <= "0000000011101000"; wait for 50 ns;
		entrada_A <= "0000000011101001"; wait for 50 ns;
		entrada_A <= "0000000011101010"; wait for 50 ns;
		entrada_A <= "0000000011101011"; wait for 50 ns;
		entrada_A <= "0000000011101100"; wait for 50 ns;
		entrada_A <= "0000000011101101"; wait for 50 ns;
		entrada_A <= "0000000011101110"; wait for 50 ns;
		entrada_A <= "0000000011101111"; wait for 50 ns;
		entrada_A <= "0000000011110000"; wait for 50 ns;
		entrada_A <= "0000000011110001"; wait for 50 ns;
		entrada_A <= "0000000011110010"; wait for 50 ns;
		entrada_A <= "0000000011110011"; wait for 50 ns;
		entrada_A <= "0000000011110100"; wait for 50 ns;
		entrada_A <= "0000000011110101"; wait for 50 ns;
		entrada_A <= "0000000011110110"; wait for 50 ns;
		entrada_A <= "0000000011110111"; wait for 50 ns;
		entrada_A <= "0000000011111000"; wait for 50 ns;
		entrada_A <= "0000000011111001"; wait for 50 ns;
		entrada_A <= "0000000011111010"; wait for 50 ns;
		entrada_A <= "0000000011111011"; wait for 50 ns;
		entrada_A <= "0000000011111100"; wait for 50 ns;
		entrada_A <= "0000000011111101"; wait for 50 ns;
		entrada_A <= "0000000011111110"; wait for 50 ns;
		entrada_A <= "0000000011111111"; wait for 50 ns;
		entrada_A <= "0000000100000000"; wait for 50 ns;
		entrada_A <= "0000000100000001"; wait for 50 ns;
		entrada_A <= "0000000100000010"; wait for 50 ns;
		entrada_A <= "0000000100000011"; wait for 50 ns;
		entrada_A <= "0000000100000100"; wait for 50 ns;
		entrada_A <= "0000000100000101"; wait for 50 ns;
		entrada_A <= "0000000100000110"; wait for 50 ns;
		entrada_A <= "0000000100000111"; wait for 50 ns;
		entrada_A <= "0000000100001000"; wait for 50 ns;
		entrada_A <= "0000000100001001"; wait for 50 ns;
		entrada_A <= "0000000100001010"; wait for 50 ns;
		entrada_A <= "0000000100001011"; wait for 50 ns;
		entrada_A <= "0000000100001100"; wait for 50 ns;
		entrada_A <= "0000000100001101"; wait for 50 ns;
		entrada_A <= "0000000100001110"; wait for 50 ns;
		entrada_A <= "0000000100001111"; wait for 50 ns;
		entrada_A <= "0000000100010000"; wait for 50 ns;
		entrada_A <= "0000000100010001"; wait for 50 ns;
		entrada_A <= "0000000100010010"; wait for 50 ns;
		entrada_A <= "0000000100010011"; wait for 50 ns;
		entrada_A <= "0000000100010100"; wait for 50 ns;
		entrada_A <= "0000000100010101"; wait for 50 ns;
		entrada_A <= "0000000100010110"; wait for 50 ns;
		entrada_A <= "0000000100010111"; wait for 50 ns;
		entrada_A <= "0000000100011000"; wait for 50 ns;
		entrada_A <= "0000000100011001"; wait for 50 ns;
		entrada_A <= "0000000100011010"; wait for 50 ns;
		entrada_A <= "0000000100011011"; wait for 50 ns;
		entrada_A <= "0000000100011100"; wait for 50 ns;
		entrada_A <= "0000000100011101"; wait for 50 ns;
		entrada_A <= "0000000100011110"; wait for 50 ns;
		entrada_A <= "0000000100011111"; wait for 50 ns;
		entrada_A <= "0000000100100000"; wait for 50 ns;
		entrada_A <= "0000000100100001"; wait for 50 ns;
		entrada_A <= "0000000100100010"; wait for 50 ns;
		entrada_A <= "0000000100100011"; wait for 50 ns;
		entrada_A <= "0000000100100100"; wait for 50 ns;
		entrada_A <= "0000000100100101"; wait for 50 ns;
		entrada_A <= "0000000100100110"; wait for 50 ns;
		entrada_A <= "0000000100100111"; wait for 50 ns;
		entrada_A <= "0000000100101000"; wait for 50 ns;
		entrada_A <= "0000000100101001"; wait for 50 ns;
		entrada_A <= "0000000100101010"; wait for 50 ns;
		entrada_A <= "0000000100101011"; wait for 50 ns;
		entrada_A <= "0000000100101100"; wait for 50 ns;
		entrada_A <= "0000000100101101"; wait for 50 ns;
		entrada_A <= "0000000100101110"; wait for 50 ns;
		entrada_A <= "0000000100101111"; wait for 50 ns;
		entrada_A <= "0000000100110000"; wait for 50 ns;
		entrada_A <= "0000000100110001"; wait for 50 ns;
		entrada_A <= "0000000100110010"; wait for 50 ns;
		entrada_A <= "0000000100110011"; wait for 50 ns;
		entrada_A <= "0000000100110100"; wait for 50 ns;
		entrada_A <= "0000000100110101"; wait for 50 ns;
		entrada_A <= "0000000100110110"; wait for 50 ns;
		entrada_A <= "0000000100110111"; wait for 50 ns;
		entrada_A <= "0000000100111000"; wait for 50 ns;
		entrada_A <= "0000000100111001"; wait for 50 ns;
		entrada_A <= "0000000100111010"; wait for 50 ns;
		entrada_A <= "0000000100111011"; wait for 50 ns;
		entrada_A <= "0000000100111100"; wait for 50 ns;
		entrada_A <= "0000000100111101"; wait for 50 ns;
		entrada_A <= "0000000100111110"; wait for 50 ns;
		entrada_A <= "0000000100111111"; wait for 50 ns;
		entrada_A <= "0000000101000000"; wait for 50 ns;
		entrada_A <= "0000000101000001"; wait for 50 ns;
		entrada_A <= "0000000101000010"; wait for 50 ns;
		entrada_A <= "0000000101000011"; wait for 50 ns;
		entrada_A <= "0000000101000100"; wait for 50 ns;
		entrada_A <= "0000000101000101"; wait for 50 ns;
		entrada_A <= "0000000101000110"; wait for 50 ns;
		entrada_A <= "0000000101000111"; wait for 50 ns;
		entrada_A <= "0000000101001000"; wait for 50 ns;
		entrada_A <= "0000000101001001"; wait for 50 ns;
		entrada_A <= "0000000101001010"; wait for 50 ns;
		entrada_A <= "0000000101001011"; wait for 50 ns;
		entrada_A <= "0000000101001100"; wait for 50 ns;
		entrada_A <= "0000000101001101"; wait for 50 ns;
		entrada_A <= "0000000101001110"; wait for 50 ns;
		entrada_A <= "0000000101001111"; wait for 50 ns;
		entrada_A <= "0000000101010000"; wait for 50 ns;
		entrada_A <= "0000000101010001"; wait for 50 ns;
		entrada_A <= "0000000101010010"; wait for 50 ns;
		entrada_A <= "0000000101010011"; wait for 50 ns;
		entrada_A <= "0000000101010100"; wait for 50 ns;
		entrada_A <= "0000000101010101"; wait for 50 ns;
		entrada_A <= "0000000101010111"; wait for 50 ns;
		entrada_A <= "0000000101011000"; wait for 50 ns;
		entrada_A <= "0000000101011001"; wait for 50 ns;
		entrada_A <= "0000000101011010"; wait for 50 ns;
		entrada_A <= "0000000101011011"; wait for 50 ns;
		entrada_A <= "0000000101011100"; wait for 50 ns;
		entrada_A <= "0000000101011101"; wait for 50 ns;
		entrada_A <= "0000000101011110"; wait for 50 ns;
		entrada_A <= "0000000101011111"; wait for 50 ns;
		entrada_A <= "0000000101100000"; wait for 50 ns;
		entrada_A <= "0000000101100001"; wait for 50 ns;
		entrada_A <= "0000000101100010"; wait for 50 ns;
		entrada_A <= "0000000101100011"; wait for 50 ns;
		entrada_A <= "0000000101100100"; wait for 50 ns;
		entrada_A <= "0000000101100101"; wait for 50 ns;
		entrada_A <= "0000000101100110"; wait for 50 ns;
		entrada_A <= "0000000101100111"; wait for 50 ns;
		entrada_A <= "0000000101101000"; wait for 50 ns;
		entrada_A <= "0000000101101001"; wait for 50 ns;
		entrada_A <= "0000000101101010"; wait for 50 ns;
		entrada_A <= "0000000101101011"; wait for 50 ns;
		entrada_A <= "0000000101101100"; wait for 50 ns;
		entrada_A <= "0000000101101101"; wait for 50 ns;
		entrada_A <= "0000000101101110"; wait for 50 ns;
		entrada_A <= "0000000101101111"; wait for 50 ns;
		entrada_A <= "0000000101110000"; wait for 50 ns;
		entrada_A <= "0000000101110001"; wait for 50 ns;
		entrada_A <= "0000000101110010"; wait for 50 ns;
		entrada_A <= "0000000101110011"; wait for 50 ns;
		entrada_A <= "0000000101110100"; wait for 50 ns;
		entrada_A <= "0000000101110101"; wait for 50 ns;
		entrada_A <= "0000000101110110"; wait for 50 ns;
		entrada_A <= "0000000101110111"; wait for 50 ns;
		entrada_A <= "0000000101111000"; wait for 50 ns;
		entrada_A <= "0000000101111001"; wait for 50 ns;
		entrada_A <= "0000000101111010"; wait for 50 ns;
		entrada_A <= "0000000101111011"; wait for 50 ns;
		entrada_A <= "0000000101111100"; wait for 50 ns;
		entrada_A <= "0000000101111101"; wait for 50 ns;
		entrada_A <= "0000000101111110"; wait for 50 ns;
		entrada_A <= "0000000101111111"; wait for 50 ns;
		entrada_A <= "0000000110000000"; wait for 50 ns;
		entrada_A <= "0000000110000001"; wait for 50 ns;
		entrada_A <= "0000000110000010"; wait for 50 ns;
		entrada_A <= "0000000110000011"; wait for 50 ns;
		entrada_A <= "0000000110000100"; wait for 50 ns;
		entrada_A <= "0000000110000101"; wait for 50 ns;
		entrada_A <= "0000000110000110"; wait for 50 ns;
		entrada_A <= "0000000110000111"; wait for 50 ns;
		entrada_A <= "0000000110001000"; wait for 50 ns;
		entrada_A <= "0000000110001001"; wait for 50 ns;
		entrada_A <= "0000000110001010"; wait for 50 ns;
		entrada_A <= "0000000110001011"; wait for 50 ns;
		entrada_A <= "0000000110001100"; wait for 50 ns;
		entrada_A <= "0000000110001101"; wait for 50 ns;
		entrada_A <= "0000000110001110"; wait for 50 ns;
		entrada_A <= "0000000110001111"; wait for 50 ns;
		entrada_A <= "0000000110010000"; wait for 50 ns;
		entrada_A <= "0000000110010001"; wait for 50 ns;
		entrada_A <= "0000000110010010"; wait for 50 ns;
		entrada_A <= "0000000110010011"; wait for 50 ns;
		entrada_A <= "0000000110010100"; wait for 50 ns;
		entrada_A <= "0000000110010101"; wait for 50 ns;
		entrada_A <= "0000000110010110"; wait for 50 ns;
		entrada_A <= "0000000110010111"; wait for 50 ns;
		entrada_A <= "0000000110011000"; wait for 50 ns;
		entrada_A <= "0000000110011001"; wait for 50 ns;
		entrada_A <= "0000000110011010"; wait for 50 ns;
		entrada_A <= "0000000110011011"; wait for 50 ns;
		entrada_A <= "0000000110011100"; wait for 50 ns;
		entrada_A <= "0000000110011101"; wait for 50 ns;
		entrada_A <= "0000000110011110"; wait for 50 ns;
		entrada_A <= "0000000110011111"; wait for 50 ns;
		entrada_A <= "0000000110100000"; wait for 50 ns;
		entrada_A <= "0000000110100001"; wait for 50 ns;
		entrada_A <= "0000000110100010"; wait for 50 ns;
		entrada_A <= "0000000110100011"; wait for 50 ns;
		entrada_A <= "0000000110100100"; wait for 50 ns;
		entrada_A <= "0000000110100101"; wait for 50 ns;
		entrada_A <= "0000000110100110"; wait for 50 ns;
		entrada_A <= "0000000110100111"; wait for 50 ns;
		entrada_A <= "0000000110101000"; wait for 50 ns;
		entrada_A <= "0000000110101001"; wait for 50 ns;
		entrada_A <= "0000000110101010"; wait for 50 ns;
		entrada_A <= "0000000110101011"; wait for 50 ns;
		entrada_A <= "0000000110101100"; wait for 50 ns;
		entrada_A <= "0000000110101101"; wait for 50 ns;
		entrada_A <= "0000000110101110"; wait for 50 ns;
		entrada_A <= "0000000110101111"; wait for 50 ns;
		entrada_A <= "0000000110110000"; wait for 50 ns;
		entrada_A <= "0000000110110001"; wait for 50 ns;
		entrada_A <= "0000000110110010"; wait for 50 ns;
		entrada_A <= "0000000110110011"; wait for 50 ns;
		entrada_A <= "0000000110110100"; wait for 50 ns;
		entrada_A <= "0000000110110101"; wait for 50 ns;
		entrada_A <= "0000000110110110"; wait for 50 ns;
		entrada_A <= "0000000110110111"; wait for 50 ns;
		entrada_A <= "0000000110111000"; wait for 50 ns;
		entrada_A <= "0000000110111001"; wait for 50 ns;
		entrada_A <= "0000000110111010"; wait for 50 ns;
		entrada_A <= "0000000110111011"; wait for 50 ns;
		entrada_A <= "0000000110111100"; wait for 50 ns;
		entrada_A <= "0000000110111101"; wait for 50 ns;
		entrada_A <= "0000000110111110"; wait for 50 ns;
		entrada_A <= "0000000110111111"; wait for 50 ns;
		entrada_A <= "0000000111000000"; wait for 50 ns;
		entrada_A <= "0000000111000001"; wait for 50 ns;
		entrada_A <= "0000000111000010"; wait for 50 ns;
		entrada_A <= "0000000111000011"; wait for 50 ns;
		entrada_A <= "0000000111000100"; wait for 50 ns;
		entrada_A <= "0000000111000101"; wait for 50 ns;
		entrada_A <= "0000000111000110"; wait for 50 ns;
		entrada_A <= "0000000111000111"; wait for 50 ns;
		entrada_A <= "0000000111001000"; wait for 50 ns;
		entrada_A <= "0000000111001001"; wait for 50 ns;
		entrada_A <= "0000000111001010"; wait for 50 ns;
		entrada_A <= "0000000111001011"; wait for 50 ns;
		entrada_A <= "0000000111001100"; wait for 50 ns;
		entrada_A <= "0000000111001101"; wait for 50 ns;
		entrada_A <= "0000000111001110"; wait for 50 ns;
		entrada_A <= "0000000111001111"; wait for 50 ns;
		entrada_A <= "0000000111010000"; wait for 50 ns;
		entrada_A <= "0000000111010001"; wait for 50 ns;
		entrada_A <= "0000000111010010"; wait for 50 ns;
		entrada_A <= "0000000111010011"; wait for 50 ns;
		entrada_A <= "0000000111010100"; wait for 50 ns;
		entrada_A <= "0000000111010101"; wait for 50 ns;
		entrada_A <= "0000000111010110"; wait for 50 ns;
		entrada_A <= "0000000111010111"; wait for 50 ns;
		entrada_A <= "0000000111011000"; wait for 50 ns;
		entrada_A <= "0000000111011001"; wait for 50 ns;
		entrada_A <= "0000000111011010"; wait for 50 ns;
		entrada_A <= "0000000111011011"; wait for 50 ns;
		entrada_A <= "0000000111011100"; wait for 50 ns;
		entrada_A <= "0000000111011101"; wait for 50 ns;
		entrada_A <= "0000000111011110"; wait for 50 ns;
		entrada_A <= "0000000111011111"; wait for 50 ns;
		entrada_A <= "0000000111100000"; wait for 50 ns;
		entrada_A <= "0000000111100001"; wait for 50 ns;
		entrada_A <= "0000000111100010"; wait for 50 ns;
		entrada_A <= "0000000111100011"; wait for 50 ns;
		entrada_A <= "0000000111100100"; wait for 50 ns;
		entrada_A <= "0000000111100101"; wait for 50 ns;
		entrada_A <= "0000000111100110"; wait for 50 ns;
		entrada_A <= "0000000111100111"; wait for 50 ns;
		entrada_A <= "0000000111101000"; wait for 50 ns;
		entrada_A <= "0000000111101001"; wait for 50 ns;
		entrada_A <= "0000000111101010"; wait for 50 ns;
		entrada_A <= "0000000111101011"; wait for 50 ns;
		entrada_A <= "0000000111101100"; wait for 50 ns;
		entrada_A <= "0000000111101101"; wait for 50 ns;
		entrada_A <= "0000000111101110"; wait for 50 ns;
		entrada_A <= "0000000111101111"; wait for 50 ns;
		entrada_A <= "0000000111110000"; wait for 50 ns;
		entrada_A <= "0000000111110001"; wait for 50 ns;
		entrada_A <= "0000000111110010"; wait for 50 ns;
		entrada_A <= "0000000111110011"; wait for 50 ns;
		entrada_A <= "0000000111110100"; wait for 50 ns;
		entrada_A <= "0000000111110101"; wait for 50 ns;
		entrada_A <= "0000000111110110"; wait for 50 ns;
		entrada_A <= "0000000111110111"; wait for 50 ns;
		entrada_A <= "0000000111111000"; wait for 50 ns;
		entrada_A <= "0000000111111001"; wait for 50 ns;
		entrada_A <= "0000000111111010"; wait for 50 ns;
		entrada_A <= "0000000111111011"; wait for 50 ns;
		entrada_A <= "0000000111111100"; wait for 50 ns;
		entrada_A <= "0000000111111101"; wait for 50 ns;
		entrada_A <= "0000000111111110"; wait for 50 ns;
		entrada_A <= "0000000111111111"; wait for 50 ns;
		entrada_A <= "0000001000000000"; wait for 50 ns;
		entrada_A <= "0000001000000001"; wait for 50 ns;
		entrada_A <= "0000001000000010"; wait for 50 ns;
		entrada_A <= "0000001000000011"; wait for 50 ns;
		entrada_A <= "0000001000000100"; wait for 50 ns;
		entrada_A <= "0000001000000101"; wait for 50 ns;
		entrada_A <= "0000001000000110"; wait for 50 ns;
		entrada_A <= "0000001000000111"; wait for 50 ns;
		entrada_A <= "0000001000001000"; wait for 50 ns;
		entrada_A <= "0000001000001001"; wait for 50 ns;
		entrada_A <= "0000001000001010"; wait for 50 ns;
		entrada_A <= "0000001000001011"; wait for 50 ns;
		entrada_A <= "0000001000001100"; wait for 50 ns;
		entrada_A <= "0000001000001101"; wait for 50 ns;
		entrada_A <= "0000001000001111"; wait for 50 ns;
		entrada_A <= "0000001000010000"; wait for 50 ns;
		entrada_A <= "0000001000010001"; wait for 50 ns;
		entrada_A <= "0000001000010010"; wait for 50 ns;
		entrada_A <= "0000001000010011"; wait for 50 ns;
		entrada_A <= "0000001000010100"; wait for 50 ns;
		entrada_A <= "0000001000010101"; wait for 50 ns;
		entrada_A <= "0000001000010110"; wait for 50 ns;
		entrada_A <= "0000001000010111"; wait for 50 ns;
		entrada_A <= "0000001000011000"; wait for 50 ns;
		entrada_A <= "0000001000011001"; wait for 50 ns;
		entrada_A <= "0000001000011010"; wait for 50 ns;
		entrada_A <= "0000001000011011"; wait for 50 ns;
		entrada_A <= "0000001000011100"; wait for 50 ns;
		entrada_A <= "0000001000011101"; wait for 50 ns;
		entrada_A <= "0000001000011110"; wait for 50 ns;
		entrada_A <= "0000001000011111"; wait for 50 ns;
		entrada_A <= "0000001000100000"; wait for 50 ns;
		entrada_A <= "0000001000100001"; wait for 50 ns;
		entrada_A <= "0000001000100010"; wait for 50 ns;
		entrada_A <= "0000001000100011"; wait for 50 ns;
		entrada_A <= "0000001000100100"; wait for 50 ns;
		entrada_A <= "0000001000100101"; wait for 50 ns;
		entrada_A <= "0000001000100110"; wait for 50 ns;
		entrada_A <= "0000001000100111"; wait for 50 ns;
		entrada_A <= "0000001000101000"; wait for 50 ns;
		entrada_A <= "0000001000101001"; wait for 50 ns;
		entrada_A <= "0000001000101010"; wait for 50 ns;
		entrada_A <= "0000001000101011"; wait for 50 ns;
		entrada_A <= "0000001000101100"; wait for 50 ns;
		entrada_A <= "0000001000101101"; wait for 50 ns;
		entrada_A <= "0000001000101110"; wait for 50 ns;
		entrada_A <= "0000001000101111"; wait for 50 ns;
		entrada_A <= "0000001000110000"; wait for 50 ns;
		entrada_A <= "0000001000110001"; wait for 50 ns;
		entrada_A <= "0000001000110010"; wait for 50 ns;
		entrada_A <= "0000001000110011"; wait for 50 ns;
		entrada_A <= "0000001000110100"; wait for 50 ns;
		entrada_A <= "0000001000110101"; wait for 50 ns;
		entrada_A <= "0000001000110110"; wait for 50 ns;
		entrada_A <= "0000001000110111"; wait for 50 ns;
		entrada_A <= "0000001000111000"; wait for 50 ns;
		entrada_A <= "0000001000111001"; wait for 50 ns;
		entrada_A <= "0000001000111010"; wait for 50 ns;
		entrada_A <= "0000001000111011"; wait for 50 ns;
		entrada_A <= "0000001000111100"; wait for 50 ns;
		entrada_A <= "0000001000111101"; wait for 50 ns;
		entrada_A <= "0000001000111110"; wait for 50 ns;
		entrada_A <= "0000001000111111"; wait for 50 ns;
		entrada_A <= "0000001001000000"; wait for 50 ns;
		entrada_A <= "0000001001000001"; wait for 50 ns;
		entrada_A <= "0000001001000010"; wait for 50 ns;
		entrada_A <= "0000001001000011"; wait for 50 ns;
		entrada_A <= "0000001001000100"; wait for 50 ns;
		entrada_A <= "0000001001000101"; wait for 50 ns;
		entrada_A <= "0000001001000110"; wait for 50 ns;
		entrada_A <= "0000001001000111"; wait for 50 ns;
		entrada_A <= "0000001001001000"; wait for 50 ns;
		entrada_A <= "0000001001001001"; wait for 50 ns;
		entrada_A <= "0000001001001010"; wait for 50 ns;
		entrada_A <= "0000001001001011"; wait for 50 ns;
		entrada_A <= "0000001001001100"; wait for 50 ns;
		entrada_A <= "0000001001001101"; wait for 50 ns;
		entrada_A <= "0000001001001110"; wait for 50 ns;
		entrada_A <= "0000001001001111"; wait for 50 ns;
		entrada_A <= "0000001001010000"; wait for 50 ns;
		entrada_A <= "0000001001010001"; wait for 50 ns;
		entrada_A <= "0000001001010010"; wait for 50 ns;
		entrada_A <= "0000001001010011"; wait for 50 ns;
		entrada_A <= "0000001001010100"; wait for 50 ns;
		entrada_A <= "0000001001010101"; wait for 50 ns;
		entrada_A <= "0000001001010110"; wait for 50 ns;
		entrada_A <= "0000001001010111"; wait for 50 ns;
		entrada_A <= "0000001001011000"; wait for 50 ns;
		entrada_A <= "0000001001011001"; wait for 50 ns;
		entrada_A <= "0000001001011010"; wait for 50 ns;
		entrada_A <= "0000001001011011"; wait for 50 ns;
		entrada_A <= "0000001001011100"; wait for 50 ns;
		entrada_A <= "0000001001011101"; wait for 50 ns;
		entrada_A <= "0000001001011110"; wait for 50 ns;
		entrada_A <= "0000001001011111"; wait for 50 ns;
		entrada_A <= "0000001001100000"; wait for 50 ns;
		entrada_A <= "0000001001100001"; wait for 50 ns;
		entrada_A <= "0000001001100010"; wait for 50 ns;
		entrada_A <= "0000001001100011"; wait for 50 ns;
		entrada_A <= "0000001001100100"; wait for 50 ns;
		entrada_A <= "0000001001100101"; wait for 50 ns;
		entrada_A <= "0000001001100110"; wait for 50 ns;
		entrada_A <= "0000001001100111"; wait for 50 ns;
		entrada_A <= "0000001001101000"; wait for 50 ns;
		entrada_A <= "0000001001101001"; wait for 50 ns;
		entrada_A <= "0000001001101010"; wait for 50 ns;
		entrada_A <= "0000001001101011"; wait for 50 ns;
		entrada_A <= "0000001001101100"; wait for 50 ns;
		entrada_A <= "0000001001101101"; wait for 50 ns;
		entrada_A <= "0000001001101110"; wait for 50 ns;
		entrada_A <= "0000001001101111"; wait for 50 ns;
		entrada_A <= "0000001001110000"; wait for 50 ns;
		entrada_A <= "0000001001110001"; wait for 50 ns;
		entrada_A <= "0000001001110010"; wait for 50 ns;
		entrada_A <= "0000001001110011"; wait for 50 ns;
		entrada_A <= "0000001001110100"; wait for 50 ns;
		entrada_A <= "0000001001110101"; wait for 50 ns;
		entrada_A <= "0000001001110110"; wait for 50 ns;
		entrada_A <= "0000001001110111"; wait for 50 ns;
		entrada_A <= "0000001001111000"; wait for 50 ns;
		entrada_A <= "0000001001111001"; wait for 50 ns;
		entrada_A <= "0000001001111010"; wait for 50 ns;
		entrada_A <= "0000001001111011"; wait for 50 ns;
		entrada_A <= "0000001001111100"; wait for 50 ns;
		entrada_A <= "0000001001111101"; wait for 50 ns;
		entrada_A <= "0000001001111110"; wait for 50 ns;
		entrada_A <= "0000001001111111"; wait for 50 ns;
		entrada_A <= "0000001010000000"; wait for 50 ns;
		entrada_A <= "0000001010000001"; wait for 50 ns;
		entrada_A <= "0000001010000010"; wait for 50 ns;
		entrada_A <= "0000001010000011"; wait for 50 ns;
		entrada_A <= "0000001010000100"; wait for 50 ns;
		entrada_A <= "0000001010000101"; wait for 50 ns;
		entrada_A <= "0000001010000110"; wait for 50 ns;
		entrada_A <= "0000001010000111"; wait for 50 ns;
		entrada_A <= "0000001010001000"; wait for 50 ns;
		entrada_A <= "0000001010001001"; wait for 50 ns;
		entrada_A <= "0000001010001010"; wait for 50 ns;
		entrada_A <= "0000001010001011"; wait for 50 ns;
		entrada_A <= "0000001010001100"; wait for 50 ns;
		entrada_A <= "0000001010001101"; wait for 50 ns;
		entrada_A <= "0000001010001110"; wait for 50 ns;
		entrada_A <= "0000001010001111"; wait for 50 ns;
		entrada_A <= "0000001010010000"; wait for 50 ns;
		entrada_A <= "0000001010010001"; wait for 50 ns;
		entrada_A <= "0000001010010010"; wait for 50 ns;
		entrada_A <= "0000001010010011"; wait for 50 ns;
		entrada_A <= "0000001010010100"; wait for 50 ns;
		entrada_A <= "0000001010010101"; wait for 50 ns;
		entrada_A <= "0000001010010110"; wait for 50 ns;
		entrada_A <= "0000001010010111"; wait for 50 ns;
		entrada_A <= "0000001010011000"; wait for 50 ns;
		entrada_A <= "0000001010011001"; wait for 50 ns;
		entrada_A <= "0000001010011010"; wait for 50 ns;
		entrada_A <= "0000001010011011"; wait for 50 ns;
		entrada_A <= "0000001010011100"; wait for 50 ns;
		entrada_A <= "0000001010011101"; wait for 50 ns;
		entrada_A <= "0000001010011110"; wait for 50 ns;
		entrada_A <= "0000001010011111"; wait for 50 ns;
		entrada_A <= "0000001010100000"; wait for 50 ns;
		entrada_A <= "0000001010100001"; wait for 50 ns;
		entrada_A <= "0000001010100010"; wait for 50 ns;
		entrada_A <= "0000001010100011"; wait for 50 ns;
		entrada_A <= "0000001010100100"; wait for 50 ns;
		entrada_A <= "0000001010100101"; wait for 50 ns;
		entrada_A <= "0000001010100110"; wait for 50 ns;
		entrada_A <= "0000001010100111"; wait for 50 ns;
		entrada_A <= "0000001010101000"; wait for 50 ns;
		entrada_A <= "0000001010010011"; wait for 50 ns;
		entrada_A <= "0000001010010100"; wait for 50 ns;
		entrada_A <= "0000001010010101"; wait for 50 ns;
		entrada_A <= "0000001010010110"; wait for 50 ns;
		entrada_A <= "0000001010010111"; wait for 50 ns;
		entrada_A <= "0000001010011000"; wait for 50 ns;
		entrada_A <= "0000001010011001"; wait for 50 ns;
		entrada_A <= "0000001010011010"; wait for 50 ns;
		entrada_A <= "0000001010011011"; wait for 50 ns;
		entrada_A <= "0000001010011100"; wait for 50 ns;
		entrada_A <= "0000001010011101"; wait for 50 ns;
		entrada_A <= "0000001010011110"; wait for 50 ns;
		entrada_A <= "0000001010011111"; wait for 50 ns;
		entrada_A <= "0000001010100000"; wait for 50 ns;
		entrada_A <= "0000001010100001"; wait for 50 ns;
		entrada_A <= "0000001010100010"; wait for 50 ns;
		entrada_A <= "0000001010100011"; wait for 50 ns;
		entrada_A <= "0000001010100100"; wait for 50 ns;
		entrada_A <= "0000001010100101"; wait for 50 ns;
		entrada_A <= "0000001010100110"; wait for 50 ns;
		entrada_A <= "0000001010100111"; wait for 50 ns;
		entrada_A <= "0000001010101000"; wait for 50 ns;
		entrada_A <= "0000001010101001"; wait for 50 ns;
		entrada_A <= "0000001010101010"; wait for 50 ns;
		entrada_A <= "0000001010101100"; wait for 50 ns;
		entrada_A <= "0000001010101101"; wait for 50 ns;
		entrada_A <= "0000001010101110"; wait for 50 ns;
		entrada_A <= "0000001010101111"; wait for 50 ns;
		entrada_A <= "0000001010110000"; wait for 50 ns;
		entrada_A <= "0000001010110001"; wait for 50 ns;
		entrada_A <= "0000001010110010"; wait for 50 ns;
		entrada_A <= "0000001010110011"; wait for 50 ns;
		entrada_A <= "0000001010110100"; wait for 50 ns;
		entrada_A <= "0000001010110101"; wait for 50 ns;
		entrada_A <= "0000001010110110"; wait for 50 ns;
		entrada_A <= "0000001010110111"; wait for 50 ns;
		entrada_A <= "0000001010111000"; wait for 50 ns;
		entrada_A <= "0000001010111001"; wait for 50 ns;
		entrada_A <= "0000001010111010"; wait for 50 ns;
		entrada_A <= "0000001010111011"; wait for 50 ns;
		entrada_A <= "0000001010111100"; wait for 50 ns;
		entrada_A <= "0000001010111101"; wait for 50 ns;
		entrada_A <= "0000001010111110"; wait for 50 ns;
		entrada_A <= "0000001010111111"; wait for 50 ns;
		entrada_A <= "0000001011000000"; wait for 50 ns;
		entrada_A <= "0000001011000001"; wait for 50 ns;
		entrada_A <= "0000001011000010"; wait for 50 ns;
		entrada_A <= "0000001011000011"; wait for 50 ns;
		entrada_A <= "0000001011000100"; wait for 50 ns;
		entrada_A <= "0000001011000101"; wait for 50 ns;
		entrada_A <= "0000001011000110"; wait for 50 ns;
		entrada_A <= "0000001011000111"; wait for 50 ns;
		entrada_A <= "0000001011001000"; wait for 50 ns;
		entrada_A <= "0000001011001001"; wait for 50 ns;
		entrada_A <= "0000001011001010"; wait for 50 ns;
		entrada_A <= "0000001011001011"; wait for 50 ns;
		entrada_A <= "0000001011001100"; wait for 50 ns;
		entrada_A <= "0000001011001101"; wait for 50 ns;
		entrada_A <= "0000001011001110"; wait for 50 ns;
		entrada_A <= "0000001011001111"; wait for 50 ns;
		entrada_A <= "0000001011010000"; wait for 50 ns;
		entrada_A <= "0000001011010001"; wait for 50 ns;
		entrada_A <= "0000001011010010"; wait for 50 ns;
		entrada_A <= "0000001011010011"; wait for 50 ns;
		entrada_A <= "0000001011010100"; wait for 50 ns;
		entrada_A <= "0000001011010101"; wait for 50 ns;
		entrada_A <= "0000001011010110"; wait for 50 ns;
		entrada_A <= "0000001011010111"; wait for 50 ns;
		entrada_A <= "0000001011011000"; wait for 50 ns;
		entrada_A <= "0000001011011001"; wait for 50 ns;
		entrada_A <= "0000001011011010"; wait for 50 ns;
		entrada_A <= "0000001011011011"; wait for 50 ns;
		entrada_A <= "0000001011011100"; wait for 50 ns;
		entrada_A <= "0000001011011101"; wait for 50 ns;
		entrada_A <= "0000001011011110"; wait for 50 ns;
		entrada_A <= "0000001011011111"; wait for 50 ns;
		entrada_A <= "0000001011100000"; wait for 50 ns;
		entrada_A <= "0000001011100001"; wait for 50 ns;
		entrada_A <= "0000001011100010"; wait for 50 ns;
		entrada_A <= "0000001011100011"; wait for 50 ns;
		entrada_A <= "0000001011100100"; wait for 50 ns;
		entrada_A <= "0000001011100101"; wait for 50 ns;
		entrada_A <= "0000001011100110"; wait for 50 ns;
		entrada_A <= "0000001011100111"; wait for 50 ns;
		entrada_A <= "0000001011101000"; wait for 50 ns;
		entrada_A <= "0000001011101001"; wait for 50 ns;
		entrada_A <= "0000001011101010"; wait for 50 ns;
		entrada_A <= "0000001011101011"; wait for 50 ns;
		entrada_A <= "0000001011101100"; wait for 50 ns;
		entrada_A <= "0000001011101101"; wait for 50 ns;
		entrada_A <= "0000001011101110"; wait for 50 ns;
		entrada_A <= "0000001011101111"; wait for 50 ns;
		entrada_A <= "0000001011110000"; wait for 50 ns;
		entrada_A <= "0000001011110001"; wait for 50 ns;
		entrada_A <= "0000001011110010"; wait for 50 ns;
		entrada_A <= "0000001011110011"; wait for 50 ns;
		entrada_A <= "0000001011110100"; wait for 50 ns;
		entrada_A <= "0000001011110101"; wait for 50 ns;
		entrada_A <= "0000001011110110"; wait for 50 ns;
		entrada_A <= "0000001011110111"; wait for 50 ns;
		entrada_A <= "0000001011111000"; wait for 50 ns;
		entrada_A <= "0000001011111001"; wait for 50 ns;
		entrada_A <= "0000001011111010"; wait for 50 ns;
		entrada_A <= "0000001011111011"; wait for 50 ns;
		entrada_A <= "0000001011111100"; wait for 50 ns;
		entrada_A <= "0000001011111101"; wait for 50 ns;
		entrada_A <= "0000001011111110"; wait for 50 ns;
		entrada_A <= "0000001011111111"; wait for 50 ns;
		entrada_A <= "0000001100000000"; wait for 50 ns;
		entrada_A <= "0000001100000001"; wait for 50 ns;
		entrada_A <= "0000001100000010"; wait for 50 ns;
		entrada_A <= "0000001100000011"; wait for 50 ns;
		entrada_A <= "0000001100000100"; wait for 50 ns;
		entrada_A <= "0000001100000101"; wait for 50 ns;
		entrada_A <= "0000001100000110"; wait for 50 ns;
		entrada_A <= "0000001100000111"; wait for 50 ns;
		entrada_A <= "0000001100001000"; wait for 50 ns;
		entrada_A <= "0000001100001001"; wait for 50 ns;
		entrada_A <= "0000001100001010"; wait for 50 ns;
		entrada_A <= "0000001100001011"; wait for 50 ns;
		entrada_A <= "0000001100001100"; wait for 50 ns;
		entrada_A <= "0000001100001101"; wait for 50 ns;
		entrada_A <= "0000001100001110"; wait for 50 ns;
		entrada_A <= "0000001100001111"; wait for 50 ns;
		entrada_A <= "0000001100010000"; wait for 50 ns;
		entrada_A <= "0000001100010001"; wait for 50 ns;
		entrada_A <= "0000001100010010"; wait for 50 ns;
		entrada_A <= "0000001100010011"; wait for 50 ns;
		entrada_A <= "0000001100010100"; wait for 50 ns;
		entrada_A <= "0000001100010101"; wait for 50 ns;
		entrada_A <= "0000001100010110"; wait for 50 ns;
		entrada_A <= "0000001100010111"; wait for 50 ns;
		entrada_A <= "0000001100011000"; wait for 50 ns;
		entrada_A <= "0000001100011001"; wait for 50 ns;
		entrada_A <= "0000001100011010"; wait for 50 ns;
		entrada_A <= "0000001100011011"; wait for 50 ns;
		entrada_A <= "0000001100011100"; wait for 50 ns;
		entrada_A <= "0000001100011101"; wait for 50 ns;
		entrada_A <= "0000001100011110"; wait for 50 ns;
		entrada_A <= "0000001100011111"; wait for 50 ns;
		entrada_A <= "0000001100100000"; wait for 50 ns;
		entrada_A <= "0000001100100001"; wait for 50 ns;
		entrada_A <= "0000001100100010"; wait for 50 ns;
		entrada_A <= "0000001100100011"; wait for 50 ns;
		entrada_A <= "0000001100100100"; wait for 50 ns;
		entrada_A <= "0000001100100101"; wait for 50 ns;
		entrada_A <= "0000001100100110"; wait for 50 ns;
		entrada_A <= "0000001100100111"; wait for 50 ns;
		entrada_A <= "0000001100101000"; wait for 50 ns;
		entrada_A <= "0000001100101001"; wait for 50 ns;
		entrada_A <= "0000001100101010"; wait for 50 ns;
		entrada_A <= "0000001100101011"; wait for 50 ns;
		entrada_A <= "0000001100101100"; wait for 50 ns;
		entrada_A <= "0000001100101101"; wait for 50 ns;
		entrada_A <= "0000001100101110"; wait for 50 ns;
		entrada_A <= "0000001100101111"; wait for 50 ns;
		entrada_A <= "0000001100110000"; wait for 50 ns;
		entrada_A <= "0000001100110001"; wait for 50 ns;
		entrada_A <= "0000001100110010"; wait for 50 ns;
		entrada_A <= "0000001100110011"; wait for 50 ns;
		entrada_A <= "0000001100110100"; wait for 50 ns;
		entrada_A <= "0000001100110101"; wait for 50 ns;
		entrada_A <= "0000001100110110"; wait for 50 ns;
		entrada_A <= "0000001100110111"; wait for 50 ns;
		entrada_A <= "0000001100111000"; wait for 50 ns;
		entrada_A <= "0000001100111001"; wait for 50 ns;
		entrada_A <= "0000001100111010"; wait for 50 ns;
		entrada_A <= "0000001100111011"; wait for 50 ns;
		entrada_A <= "0000001100111100"; wait for 50 ns;
		entrada_A <= "0000001100111101"; wait for 50 ns;
		entrada_A <= "0000001100111110"; wait for 50 ns;
		entrada_A <= "0000001100111111"; wait for 50 ns;
		entrada_A <= "0000001101000000"; wait for 50 ns;
		entrada_A <= "0000001101000001"; wait for 50 ns;
		entrada_A <= "0000001101000010"; wait for 50 ns;
		entrada_A <= "0000001101000011"; wait for 50 ns;
		entrada_A <= "0000001101000100"; wait for 50 ns;
		entrada_A <= "0000001101000101"; wait for 50 ns;
		entrada_A <= "0000001101000110"; wait for 50 ns;
		entrada_A <= "0000001101000111"; wait for 50 ns;
		entrada_A <= "0000001101001000"; wait for 50 ns;
		entrada_A <= "0000001101001001"; wait for 50 ns;
		entrada_A <= "0000001101001010"; wait for 50 ns;
		entrada_A <= "0000001101001011"; wait for 50 ns;
		entrada_A <= "0000001101001100"; wait for 50 ns;
		entrada_A <= "0000001101001101"; wait for 50 ns;
		entrada_A <= "0000001101001110"; wait for 50 ns;
		entrada_A <= "0000001101001111"; wait for 50 ns;
		entrada_A <= "0000001101010000"; wait for 50 ns;
		entrada_A <= "0000001101010001"; wait for 50 ns;
		entrada_A <= "0000001101010010"; wait for 50 ns;
		entrada_A <= "0000001101010011"; wait for 50 ns;
		entrada_A <= "0000001101010100"; wait for 50 ns;
		entrada_A <= "0000001101010101"; wait for 50 ns;
		entrada_A <= "0000001101010111"; wait for 50 ns;
		entrada_A <= "0000001101011000"; wait for 50 ns;
		entrada_A <= "0000001101011001"; wait for 50 ns;
		entrada_A <= "0000001101011010"; wait for 50 ns;
		entrada_A <= "0000001101011011"; wait for 50 ns;
		entrada_A <= "0000001101011100"; wait for 50 ns;
		entrada_A <= "0000001101011101"; wait for 50 ns;
		entrada_A <= "0000001101011110"; wait for 50 ns;
		entrada_A <= "0000001101011111"; wait for 50 ns;
		entrada_A <= "0000001101100000"; wait for 50 ns;
		entrada_A <= "0000001101100001"; wait for 50 ns;
		entrada_A <= "0000001101100010"; wait for 50 ns;
		entrada_A <= "0000001101100011"; wait for 50 ns;
		entrada_A <= "0000001101100100"; wait for 50 ns;
		entrada_A <= "0000001101100101"; wait for 50 ns;
		entrada_A <= "0000001101100110"; wait for 50 ns;
		entrada_A <= "0000001101100111"; wait for 50 ns;
		entrada_A <= "0000001101101000"; wait for 50 ns;
		entrada_A <= "0000001101101001"; wait for 50 ns;
		entrada_A <= "0000001101101010"; wait for 50 ns;
		entrada_A <= "0000001101101011"; wait for 50 ns;
		entrada_A <= "0000001101101100"; wait for 50 ns;
		entrada_A <= "0000001101101101"; wait for 50 ns;
		entrada_A <= "0000001101101110"; wait for 50 ns;
		entrada_A <= "0000001101101111"; wait for 50 ns;
		entrada_A <= "0000001101110000"; wait for 50 ns;
		entrada_A <= "0000001101110001"; wait for 50 ns;
		entrada_A <= "0000001101110010"; wait for 50 ns;
		entrada_A <= "0000001101110011"; wait for 50 ns;
		entrada_A <= "0000001101110100"; wait for 50 ns;
		entrada_A <= "0000001101110101"; wait for 50 ns;
		entrada_A <= "0000001101110110"; wait for 50 ns;
		entrada_A <= "0000001101110111"; wait for 50 ns;
		entrada_A <= "0000001101111000"; wait for 50 ns;
		entrada_A <= "0000001101111001"; wait for 50 ns;
		entrada_A <= "0000001101111010"; wait for 50 ns;
		entrada_A <= "0000001101111011"; wait for 50 ns;
		entrada_A <= "0000001101111100"; wait for 50 ns;
		entrada_A <= "0000001101111101"; wait for 50 ns;
		entrada_A <= "0000001101111110"; wait for 50 ns;
		entrada_A <= "0000001101111111"; wait for 50 ns;
		entrada_A <= "0000001110000000"; wait for 50 ns;
		entrada_A <= "0000001110000001"; wait for 50 ns;
		entrada_A <= "0000001110000010"; wait for 50 ns;
		entrada_A <= "0000001110000011"; wait for 50 ns;
		entrada_A <= "0000001110000100"; wait for 50 ns;
		entrada_A <= "0000001110000101"; wait for 50 ns;
		entrada_A <= "0000001110000110"; wait for 50 ns;
		entrada_A <= "0000001110000111"; wait for 50 ns;
		entrada_A <= "0000001110001000"; wait for 50 ns;
		entrada_A <= "0000001110001001"; wait for 50 ns;
		entrada_A <= "0000001110001010"; wait for 50 ns;
		entrada_A <= "0000001110001011"; wait for 50 ns;
		entrada_A <= "0000001110001100"; wait for 50 ns;
		entrada_A <= "0000001110001101"; wait for 50 ns;
		entrada_A <= "0000001110001110"; wait for 50 ns;
		entrada_A <= "0000001110001111"; wait for 50 ns;
		entrada_A <= "0000001110010000"; wait for 50 ns;
		entrada_A <= "0000001110010001"; wait for 50 ns;
		entrada_A <= "0000001110010010"; wait for 50 ns;
		entrada_A <= "0000001110010011"; wait for 50 ns;
		entrada_A <= "0000001110010100"; wait for 50 ns;
		entrada_A <= "0000001110010101"; wait for 50 ns;
		entrada_A <= "0000001110010110"; wait for 50 ns;
		entrada_A <= "0000001110010111"; wait for 50 ns;
		entrada_A <= "0000001110011000"; wait for 50 ns;
		entrada_A <= "0000001110011001"; wait for 50 ns;
		entrada_A <= "0000001110011010"; wait for 50 ns;
		entrada_A <= "0000001110011011"; wait for 50 ns;
		entrada_A <= "0000001110011100"; wait for 50 ns;
		entrada_A <= "0000001110011101"; wait for 50 ns;
		entrada_A <= "0000001110011110"; wait for 50 ns;
		entrada_A <= "0000001110011111"; wait for 50 ns;
		entrada_A <= "0000001110100000"; wait for 50 ns;
		entrada_A <= "0000001110100001"; wait for 50 ns;
		entrada_A <= "0000001110100010"; wait for 50 ns;
		entrada_A <= "0000001110100011"; wait for 50 ns;
		entrada_A <= "0000001110100100"; wait for 50 ns;
		entrada_A <= "0000001110100101"; wait for 50 ns;
		entrada_A <= "0000001110100110"; wait for 50 ns;
		entrada_A <= "0000001110100111"; wait for 50 ns;
		entrada_A <= "0000001110101000"; wait for 50 ns;
		entrada_A <= "0000001110101001"; wait for 50 ns;
		entrada_A <= "0000001110101010"; wait for 50 ns;
		entrada_A <= "0000001110101011"; wait for 50 ns;
		entrada_A <= "0000001110101100"; wait for 50 ns;
		entrada_A <= "0000001110101101"; wait for 50 ns;
		entrada_A <= "0000001110101110"; wait for 50 ns;
		entrada_A <= "0000001110101111"; wait for 50 ns;
		entrada_A <= "0000001110110000"; wait for 50 ns;
		entrada_A <= "0000001110110001"; wait for 50 ns;
		entrada_A <= "0000001110110010"; wait for 50 ns;
		entrada_A <= "0000001110110011"; wait for 50 ns;
		entrada_A <= "0000001110110100"; wait for 50 ns;
		entrada_A <= "0000001110110101"; wait for 50 ns;
		entrada_A <= "0000001110110110"; wait for 50 ns;
		entrada_A <= "0000001110110111"; wait for 50 ns;
		entrada_A <= "0000001110111000"; wait for 50 ns;
		entrada_A <= "0000001110111001"; wait for 50 ns;
		entrada_A <= "0000001110111010"; wait for 50 ns;
		entrada_A <= "0000001110111011"; wait for 50 ns;
		entrada_A <= "0000001110111100"; wait for 50 ns;
		entrada_A <= "0000001110111101"; wait for 50 ns;
		entrada_A <= "0000001110111110"; wait for 50 ns;
		entrada_A <= "0000001110111111"; wait for 50 ns;
		entrada_A <= "0000001111000000"; wait for 50 ns;
		entrada_A <= "0000001111000001"; wait for 50 ns;
		entrada_A <= "0000001111000010"; wait for 50 ns;
		entrada_A <= "0000001111000011"; wait for 50 ns;
		entrada_A <= "0000001111000100"; wait for 50 ns;
		entrada_A <= "0000001111000101"; wait for 50 ns;
		entrada_A <= "0000001111000110"; wait for 50 ns;
		entrada_A <= "0000001111000111"; wait for 50 ns;
		entrada_A <= "0000001111001000"; wait for 50 ns;
		entrada_A <= "0000001111001001"; wait for 50 ns;
		entrada_A <= "0000001111001010"; wait for 50 ns;
		entrada_A <= "0000001111001011"; wait for 50 ns;
		entrada_A <= "0000001111001100"; wait for 50 ns;
		entrada_A <= "0000001111001101"; wait for 50 ns;
		entrada_A <= "0000001111001110"; wait for 50 ns;
		entrada_A <= "0000001111001111"; wait for 50 ns;
		entrada_A <= "0000001111010000"; wait for 50 ns;
		entrada_A <= "0000001111010001"; wait for 50 ns;
		entrada_A <= "0000001111010010"; wait for 50 ns;
		entrada_A <= "0000001111010011"; wait for 50 ns;
		entrada_A <= "0000001111010100"; wait for 50 ns;
		entrada_A <= "0000001111010101"; wait for 50 ns;
		entrada_A <= "0000001111010110"; wait for 50 ns;
		entrada_A <= "0000001111010111"; wait for 50 ns;
		entrada_A <= "0000001111011000"; wait for 50 ns;
		entrada_A <= "0000001111011001"; wait for 50 ns;
		entrada_A <= "0000001111011010"; wait for 50 ns;
		entrada_A <= "0000001111011011"; wait for 50 ns;
		entrada_A <= "0000001111011100"; wait for 50 ns;
		entrada_A <= "0000001111011101"; wait for 50 ns;
		entrada_A <= "0000001111011110"; wait for 50 ns;
		entrada_A <= "0000001111011111"; wait for 50 ns;
		entrada_A <= "0000001111100000"; wait for 50 ns;
		entrada_A <= "0000001111100001"; wait for 50 ns;
		entrada_A <= "0000001111100010"; wait for 50 ns;
		entrada_A <= "0000001111100011"; wait for 50 ns;
		entrada_A <= "0000001111100100"; wait for 50 ns;
		entrada_A <= "0000001111100101"; wait for 50 ns;
		entrada_A <= "0000001111100110"; wait for 50 ns;
		entrada_A <= "0000001111100111"; wait for 50 ns;
		entrada_A <= "0000001111101000"; wait for 50 ns;
		entrada_A <= "0000001111101001"; wait for 50 ns;
		entrada_A <= "0000001111101010"; wait for 50 ns;
		entrada_A <= "0000001111101011"; wait for 50 ns;
		entrada_A <= "0000001111101100"; wait for 50 ns;
		entrada_A <= "0000001111101101"; wait for 50 ns;
		entrada_A <= "0000001111101110"; wait for 50 ns;
		entrada_A <= "0000001111101111"; wait for 50 ns;
		entrada_A <= "0000001111110000"; wait for 50 ns;
		entrada_A <= "0000001111110001"; wait for 50 ns;
		entrada_A <= "0000001111110010"; wait for 50 ns;
		entrada_A <= "0000001111110011"; wait for 50 ns;
		entrada_A <= "0000001111110100"; wait for 50 ns;
		entrada_A <= "0000001111110101"; wait for 50 ns;
		entrada_A <= "0000001111110110"; wait for 50 ns;
		entrada_A <= "0000001111110111"; wait for 50 ns;
		entrada_A <= "0000001111111000"; wait for 50 ns;
		entrada_A <= "0000001111111001"; wait for 50 ns;
		entrada_A <= "0000001111111010"; wait for 50 ns;
		entrada_A <= "0000001111111011"; wait for 50 ns;
		entrada_A <= "0000001111111100"; wait for 50 ns;
		entrada_A <= "0000001111111101"; wait for 50 ns;
		entrada_A <= "0000001111111110"; wait for 50 ns;
		entrada_A <= "0000001111111111"; wait for 50 ns;
		entrada_A <= "0000010000000000"; wait for 50 ns;
	end process;
	
	signal_b_somador : process
	begin
	
	end process;
end hardware;